
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_omp_reconstruction.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_omp_reconstruction.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_omp_reconstruction.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = 1'b0;
    assign module_intf_7.ap_ready = 1'b0;
    assign module_intf_7.ap_done = 1'b0;
    assign module_intf_7.ap_continue = 1'b0;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = 1'b0;
    assign module_intf_10.ap_ready = 1'b0;
    assign module_intf_10.ap_done = 1'b0;
    assign module_intf_10.ap_continue = 1'b0;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;

    seq_loop_intf#(182) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state9;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state13;
    assign seq_loop_intf_1.post_states_valid = 1'b1;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state10;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_omp_reconstruction.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_omp_reconstruction.ap_ST_fsm_state10;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state12;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(182) seq_loop_monitor_1;
    seq_loop_intf#(182) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state14;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state17;
    assign seq_loop_intf_2.post_states_valid = 1'b1;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state15;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_omp_reconstruction.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_omp_reconstruction.ap_ST_fsm_state15;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state16;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(182) seq_loop_monitor_2;
    seq_loop_intf#(182) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state17;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state20;
    assign seq_loop_intf_3.post_states_valid = 1'b1;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state18;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_omp_reconstruction.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_omp_reconstruction.ap_ST_fsm_state18;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state19;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(182) seq_loop_monitor_3;
    seq_loop_intf#(182) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state10;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state122;
    assign seq_loop_intf_4.post_states_valid = 1'b1;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state13;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_omp_reconstruction.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_omp_reconstruction.ap_ST_fsm_state13;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_omp_reconstruction.ap_ST_fsm_state121;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(182) seq_loop_monitor_4;
    seq_loop_intf#(220) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state3;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state6;
    assign seq_loop_intf_5.post_states_valid = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state4;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state4;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state5;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(220) seq_loop_monitor_5;
    seq_loop_intf#(220) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state1;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state108;
    assign seq_loop_intf_6.post_states_valid = 1'b1;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state2;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state2;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_omp_reconstruction.grp_gram_schmidt_fu_3826.ap_ST_fsm_state107;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(220) seq_loop_monitor_6;
    seq_loop_intf#(134) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state33;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state41;
    assign seq_loop_intf_7.post_states_valid = 1'b1;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state34;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state34;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state40;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(134) seq_loop_monitor_7;
    seq_loop_intf#(134) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state47;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state55;
    assign seq_loop_intf_8.post_states_valid = 1'b1;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state48;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state48;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state54;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(134) seq_loop_monitor_8;
    seq_loop_intf#(134) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state61;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state69;
    assign seq_loop_intf_9.post_states_valid = 1'b1;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state62;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state62;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state68;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(134) seq_loop_monitor_9;
    seq_loop_intf#(134) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state75;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state83;
    assign seq_loop_intf_10.post_states_valid = 1'b1;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state76;
    assign seq_loop_intf_10.quit_states_valid = 1'b1;
    assign seq_loop_intf_10.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state76;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state82;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(134) seq_loop_monitor_10;
    seq_loop_intf#(134) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state89;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state97;
    assign seq_loop_intf_11.post_states_valid = 1'b1;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state90;
    assign seq_loop_intf_11.quit_states_valid = 1'b1;
    assign seq_loop_intf_11.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state90;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state96;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(134) seq_loop_monitor_11;
    seq_loop_intf#(134) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state103;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state111;
    assign seq_loop_intf_12.post_states_valid = 1'b1;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state104;
    assign seq_loop_intf_12.quit_states_valid = 1'b1;
    assign seq_loop_intf_12.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state104;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state110;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(134) seq_loop_monitor_12;
    seq_loop_intf#(134) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state6;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state118;
    assign seq_loop_intf_13.post_states_valid = 1'b1;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state7;
    assign seq_loop_intf_13.quit_states_valid = 1'b1;
    assign seq_loop_intf_13.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state7;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state117;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(134) seq_loop_monitor_13;
    seq_loop_intf#(134) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state122;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state121;
    assign seq_loop_intf_14.post_states_valid = 1'b1;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state123;
    assign seq_loop_intf_14.quit_states_valid = 1'b1;
    assign seq_loop_intf_14.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state123;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state127;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(134) seq_loop_monitor_14;
    seq_loop_intf#(134) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state120;
    assign seq_loop_intf_15.pre_states_valid = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state120;
    assign seq_loop_intf_15.post_states_valid = 1'b1;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state121;
    assign seq_loop_intf_15.quit_states_valid = 1'b1;
    assign seq_loop_intf_15.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state121;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state123;
    assign seq_loop_intf_15.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(134) seq_loop_monitor_15;
    seq_loop_intf#(134) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state119;
    assign seq_loop_intf_16.pre_states_valid = 1'b1;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state128;
    assign seq_loop_intf_16.post_states_valid = 1'b1;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state120;
    assign seq_loop_intf_16.quit_states_valid = 1'b1;
    assign seq_loop_intf_16.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state120;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.ap_ST_fsm_state121;
    assign seq_loop_intf_16.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(134) seq_loop_monitor_16;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_init_x_fu_3663.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_2.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_load_A_col_fu_3670.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_enable_reg_pp0_iter100;
    assign upc_loop_intf_3.quit_enable = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_enable_reg_pp0_iter100;
    assign upc_loop_intf_3.loop_start = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_omp_reconstruction.grp_atom_selection_fu_3726.grp_atom_selection_Pipeline_atom_loop_fu_1118.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_enable_reg_pp0_iter99;
    assign upc_loop_intf_4.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_enable_reg_pp0_iter99;
    assign upc_loop_intf_4.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_G_VITIS_LOOP_254_1_fu_4027.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_enable_reg_pp0_iter99;
    assign upc_loop_intf_5.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_enable_reg_pp0_iter99;
    assign upc_loop_intf_5.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_compute_b_fu_4087.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(1) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1;
    assign upc_loop_intf_6.quit_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_6.quit_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_6.iter_start_enable = 1'b1;
    assign upc_loop_intf_6.iter_end_enable = 1'b1;
    assign upc_loop_intf_6.quit_enable = 1'b1;
    assign upc_loop_intf_6.loop_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_init_mats_fu_2762.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b1;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(1) upc_loop_monitor_6;
    upc_loop_intf#(1) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_7.quit_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_enable_reg_pp0_iter5;
    assign upc_loop_intf_7.loop_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_inv_d_loop_fu_2886.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(1) upc_loop_monitor_7;
    upc_loop_intf#(1) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.loop_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_T_fu_2906.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(1) upc_loop_monitor_8;
    upc_loop_intf#(1) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_9.quit_enable = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_enable_reg_pp0_iter18;
    assign upc_loop_intf_9.loop_start = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_omp_reconstruction.grp_acd_inversion_fu_4195.grp_acd_inversion_Pipeline_calc_Ginv_fu_3060.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(1) upc_loop_monitor_9;
    upc_loop_intf#(1) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_10.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_enable_reg_pp0_iter17;
    assign upc_loop_intf_10.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_mult_theta_fu_4273.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b1;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(1) upc_loop_monitor_10;
    upc_loop_intf#(1) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_enable_reg_pp0_iter8;
    assign upc_loop_intf_11.quit_enable = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_enable_reg_pp0_iter8;
    assign upc_loop_intf_11.loop_start = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_omp_reconstruction.grp_omp_reconstruction_Pipeline_map_out_fu_4350.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b1;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(1) upc_loop_monitor_11;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
